`timescale 1ns/1ns;
module shifter_tb();
    reg [15:0]  shift_in;
    reg [3:0]   shift_val;
    reg [1:0]   mode;
    wire [15:0] shift_out;
    wire [2:0]  flag;

    initial begin
    end

    initial begin
    end

endmodule