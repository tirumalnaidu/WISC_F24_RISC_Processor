`ifndef _FLAGS_H
`define _FLAGS_H
`define FLAG_Z 0
`define FLAG_V 1
`define FLAG_N 2
`endif